ibrary IEEE;
use IEEE.std_logic_1164.all;
use std.textio.all;

entity test3_tb is
end test3_tb;

architecture a_test3_tb of test3_tb is

constant C_FILE_NAME :string  := "DataOut.dat";

component test3 is
