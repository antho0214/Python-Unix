Library IEEE;
use IEEE.std_logic_1164.all;
use std.textio.all;
entity mul8u_17C8 is
port (A : in std_logic_vector(7 downto 0);
B : in std_logic_vector(7 downto 0);
O : out std_logic_vector(15 downto 0)
);
end mul8u_17C8;
architecture mul8u_17C8_struct of mul8u_17C8 is
signal sig_52,sig_53,sig_85,sig_95,sig_96,sig_127,sig_128,sig_130,sig_137,sig_138,sig_139,sig_165,sig_166,sig_170,sig_171,sig_173,sig_174,sig_180,sig_181,sig_182: std_logic;
signal sig_199,sig_208,sig_209,sig_210,sig_211,sig_212,sig_213,sig_214,sig_215,sig_216,sig_217,sig_222,sig_223,sig_224,sig_225,sig_239,sig_246,sig_247,sig_248,sig_249: std_logic;
signal sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256,sig_257,sig_258,sig_259,sig_260,sig_263,sig_264,sig_265,sig_266,sig_267,sig_268,sig_284,sig_285,sig_286: std_logic;
signal sig_287,sig_288,sig_289,sig_290,sig_291,sig_292,sig_293,sig_294,sig_295,sig_296,sig_297,sig_298,sig_299,sig_300,sig_301,sig_302,sig_303,sig_309,sig_313,sig_316: std_logic;
signal sig_317,sig_318,sig_319,sig_320,sig_321,sig_322,sig_323,sig_324,sig_325,sig_326,sig_327,sig_328,sig_329,sig_330,sig_331,sig_332,sig_333,sig_334,sig_335: std_logic;
begin
sig_52 <= B(7) and A(2);
sig_53 <= B(7) and A(2);
sig_85 <= A(3) and sig_52;
sig_95 <= B(6) and A(3);
sig_96 <= B(7) and A(3);
sig_127 <= sig_53 xor sig_95;
sig_128 <= sig_53 and A(3);
sig_130 <= sig_127 xor sig_85;
sig_137 <= B(5) and A(4);
sig_138 <= B(6) and A(4);
sig_139 <= B(7) and A(4);
sig_165 <= sig_130 or sig_137;
sig_166 <= sig_130 and sig_137;
sig_170 <= sig_96 xor sig_138;
sig_171 <= sig_96 and sig_138;
sig_173 <= sig_170 xor sig_85;
sig_174 <= sig_171 or sig_128;
sig_180 <= B(5) and A(5);
sig_181 <= B(6) and A(5);
sig_182 <= B(7) and A(5);
sig_199 <= B(3) and A(6);
sig_208 <= sig_173 xor sig_180;
sig_209 <= sig_173 and sig_180;
sig_210 <= sig_208 and sig_166;
sig_211 <= sig_208 xor sig_166;
sig_212 <= sig_209 or sig_210;
sig_213 <= sig_139 xor sig_181;
sig_214 <= sig_139 and sig_181;
sig_215 <= sig_213 and sig_174;
sig_216 <= sig_213 xor sig_174;
sig_217 <= sig_214 or sig_215;
sig_222 <= B(4) and A(6);
sig_223 <= B(5) and A(6);
sig_224 <= B(6) and A(6);
sig_225 <= B(7) and A(6);
sig_239 <= A(5) and B(4);
sig_246 <= sig_211 xor sig_222;
sig_247 <= sig_211 and sig_222;
sig_248 <= sig_246 and sig_165;
sig_249 <= sig_246 xor sig_165;
sig_250 <= sig_247 or sig_248;
sig_251 <= sig_216 xor sig_223;
sig_252 <= sig_216 and sig_223;
sig_253 <= sig_251 and sig_212;
sig_254 <= sig_251 xor sig_212;
sig_255 <= sig_252 or sig_253;
sig_256 <= sig_182 xor sig_224;
sig_257 <= sig_182 and sig_224;
sig_258 <= sig_256 and sig_217;
sig_259 <= sig_256 xor sig_217;
sig_260 <= sig_257 or sig_258;
sig_263 <= B(2) and A(7);
sig_264 <= B(3) and A(7);
sig_265 <= B(4) and A(7);
sig_266 <= B(5) and A(7);
sig_267 <= B(6) and A(7);
sig_268 <= B(7) and A(7);
sig_284 <= sig_249 xor sig_264;
sig_285 <= sig_249 and sig_264;
sig_286 <= sig_284 and sig_199;
sig_287 <= sig_284 xor sig_199;
sig_288 <= sig_285 or sig_286;
sig_289 <= sig_254 xor sig_265;
sig_290 <= sig_254 and sig_265;
sig_291 <= sig_289 and sig_250;
sig_292 <= sig_289 xor sig_250;
sig_293 <= sig_290 or sig_291;
sig_294 <= sig_259 xor sig_266;
sig_295 <= sig_259 and sig_266;
sig_296 <= sig_294 and sig_255;
sig_297 <= sig_294 xor sig_255;
sig_298 <= sig_295 or sig_296;
sig_299 <= sig_225 xor sig_267;
sig_300 <= sig_225 and sig_267;
sig_301 <= sig_299 and sig_260;
sig_302 <= sig_299 xor sig_260;
sig_303 <= sig_300 or sig_301;
sig_309 <= sig_239 xor sig_263;
sig_313 <= sig_239 and sig_263;
sig_316 <= sig_292 xor sig_288;
sig_317 <= sig_292 and sig_288;
sig_318 <= sig_316 and sig_313;
sig_319 <= sig_316 xor sig_313;
sig_320 <= sig_317 or sig_318;
sig_321 <= sig_297 xor sig_293;
sig_322 <= sig_297 and sig_293;
sig_323 <= sig_321 and sig_320;
sig_324 <= sig_321 xor sig_320;
sig_325 <= sig_322 or sig_323;
sig_326 <= sig_302 xor sig_298;
sig_327 <= sig_302 and sig_298;
sig_328 <= sig_326 and sig_325;
sig_329 <= sig_326 xor sig_325;
sig_330 <= sig_327 or sig_328;
sig_331 <= sig_268 xor sig_303;
sig_332 <= A(7) and sig_303;
sig_333 <= sig_268 and sig_330;
sig_334 <= sig_331 xor sig_330;
sig_335 <= sig_332 or sig_333;
O(15) <= sig_335;
O(14) <= sig_334;
O(13) <= sig_329;
O(12) <= sig_324;
O(11) <= sig_319;
O(10) <= sig_287;
O(9) <= sig_309;
O(8) <= sig_309;
O(7) <= sig_214;
O(6) <= sig_254;
O(5) <= sig_225;
O(4) <= sig_127;
O(3) <= '0';
O(2) <= sig_309;
O(1) <= sig_291;
O(0) <= sig_217;
end mul8u_17C8_struct;
