Library IEEE;
use IEEE.std_logic_1164.all;
use std.textio.all;
entity mul8u_T83 is
port (A : in std_logic_vector(7 downto 0);
B : in std_logic_vector(7 downto 0);
O : out std_logic_vector(15 downto 0)
);
end mul8u_T83;
architecture mul8u_T83_struct of mul8u_T83 is
signal sig_138,sig_139,sig_171,sig_181,sig_182,sig_209,sig_213,sig_216,sig_224,sig_225,sig_247,sig_256,sig_257,sig_259,sig_265,sig_266,sig_267,sig_268,sig_293,sig_294: std_logic;
signal sig_295,sig_296,sig_297,sig_298,sig_299,sig_300,sig_301,sig_302,sig_303,sig_321,sig_322,sig_323,sig_324,sig_325,sig_326,sig_327,sig_328,sig_329,sig_330,sig_331: std_logic;
signal sig_332: std_logic;
begin
sig_138 <= B(6) and A(5);
sig_139 <= B(7) and A(4);
sig_171 <= B(7) and sig_138;
sig_181 <= B(6) and A(5);
sig_182 <= B(7) and A(5);
sig_209 <= A(6) and B(5);
sig_213 <= sig_139 xor sig_181;
sig_216 <= sig_213 xor sig_171;
sig_224 <= B(6) and A(6);
sig_225 <= B(7) and A(6);
sig_247 <= B(3) and A(3);
sig_256 <= sig_182 xor sig_224;
sig_257 <= sig_182 and sig_181;
sig_259 <= sig_256 xor sig_171;
sig_265 <= B(4) and A(7);
sig_266 <= B(5) and A(7);
sig_267 <= B(6) and A(7);
sig_268 <= B(7) and A(7);
sig_293 <= sig_265 or sig_247;
sig_294 <= sig_259 xor sig_266;
sig_295 <= sig_259 and sig_266;
sig_296 <= sig_294 and sig_209;
sig_297 <= sig_294 xor sig_209;
sig_298 <= sig_295 or sig_296;
sig_299 <= sig_225 xor sig_267;
sig_300 <= sig_225 and sig_267;
sig_301 <= sig_299 and sig_257;
sig_302 <= sig_299 xor sig_257;
sig_303 <= sig_300 or sig_301;
sig_321 <= sig_297 xor sig_293;
sig_322 <= sig_297 and sig_293;
sig_323 <= sig_302 xor sig_298;
sig_324 <= sig_302 and sig_298;
sig_325 <= sig_323 and sig_322;
sig_326 <= sig_323 xor sig_322;
sig_327 <= sig_324 or sig_325;
sig_328 <= sig_268 xor sig_303;
sig_329 <= A(7) and sig_303;
sig_330 <= sig_268 and sig_327;
sig_331 <= sig_328 xor sig_327;
sig_332 <= sig_329 or sig_330;
O(15) <= sig_332;
O(14) <= sig_331;
O(13) <= sig_326;
O(12) <= sig_321;
O(11) <= sig_216;
O(10) <= sig_216;
O(9) <= sig_321;
O(8) <= sig_216;
O(7) <= sig_139;
O(6) <= sig_181;
O(5) <= sig_303;
O(4) <= '0';
O(3) <= '0';
O(2) <= sig_326;
O(1) <= '0';
O(0) <= '0';
end mul8u_T83_struct;
