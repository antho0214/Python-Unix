entity mul8u_197B is
port (A : in std_logic_vector (7 downto 0);
B : in std_logic_vector (7 downto 0);
O : out std_logic_vector (15 downto 0)
);
end mul8u_197B;
architecture mul8u_197B_struct of mul8u_197B is
signal sig_23,sig_24,sig_30,sig_31,sig_44,sig_45,sig_52,sig_53,sig_79,sig_80,sig_82,sig_85,sig_87,sig_88,sig_93,sig_94,sig_95,sig_96,sig_113,sig_117: std_logic;
signal sig_118,sig_122,sig_123,sig_124,sig_125,sig_126,sig_127,sig_128,sig_129,sig_130,sig_131,sig_136,sig_137,sig_138,sig_139,sig_160,sig_161,sig_162,sig_163,sig_164: std_logic;
signal sig_165,sig_166,sig_167,sig_168,sig_169,sig_170,sig_171,sig_172,sig_173,sig_174,sig_177,sig_178,sig_179,sig_180,sig_181,sig_182,sig_196,sig_198,sig_199,sig_200: std_logic;
signal sig_201,sig_202,sig_203,sig_204,sig_205,sig_206,sig_207,sig_208,sig_209,sig_210,sig_211,sig_212,sig_213,sig_214,sig_215,sig_216,sig_217,sig_219,sig_220,sig_221: std_logic;
signal sig_222,sig_223,sig_224,sig_225,sig_231,sig_232,sig_236,sig_237,sig_238,sig_239,sig_240,sig_241,sig_242,sig_243,sig_244,sig_245,sig_246,sig_247,sig_248,sig_249: std_logic;
signal sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256,sig_257,sig_258,sig_259,sig_260,sig_261,sig_262,sig_263,sig_264,sig_265,sig_266,sig_267,sig_268,sig_273: std_logic;
signal sig_274,sig_275,sig_276,sig_277,sig_278,sig_279,sig_280,sig_281,sig_282,sig_283,sig_284,sig_285,sig_286,sig_287,sig_288,sig_289,sig_290,sig_291,sig_292,sig_293: std_logic;
signal sig_294,sig_295,sig_296,sig_297,sig_298,sig_299,sig_301,sig_302,sig_303,sig_306,sig_307,sig_311,sig_312,sig_313,sig_314,sig_315,sig_316,sig_317,sig_318,sig_319: std_logic;
signal sig_320,sig_321,sig_322,sig_323,sig_324,sig_325,sig_326,sig_327,sig_328,sig_329,sig_330,sig_331,sig_332,sig_333,sig_334,sig_335: std_logic;
begin
sig_23 <= B(7) and A(0);
sig_24 <= A(2) and B(5);
sig_30 <= B(6) and A(1);
sig_31 <= B(7) and A(1);
sig_44 <= sig_23 or sig_30;
sig_45 <= sig_23 and sig_30;
sig_52 <= B(6) and A(2);
sig_53 <= B(7) and A(2);
sig_79 <= sig_44 xor A(4);
sig_80 <= sig_52 xor sig_31;
sig_82 <= sig_79 xor A(4);
sig_85 <= sig_31 and sig_52;
sig_87 <= sig_80 xor sig_45;
sig_88 <= sig_85 or sig_45;
sig_93 <= B(4) and A(3);
sig_94 <= B(5) and A(3);
sig_95 <= B(6) and A(3);
sig_96 <= B(7) and A(3);
sig_113 <= B(3) and A(4);
sig_117 <= sig_82 or sig_93;
sig_118 <= sig_82 and sig_93;
sig_122 <= sig_87 xor sig_94;
sig_123 <= sig_87 and sig_94;
sig_124 <= sig_122 and sig_24;
sig_125 <= sig_122 xor sig_24;
sig_126 <= sig_123 or sig_124;
sig_127 <= sig_53 xor sig_95;
sig_128 <= sig_53 and sig_95;
sig_129 <= sig_127 and sig_88;
sig_130 <= sig_127 xor sig_88;
sig_131 <= sig_128 or sig_129;
sig_136 <= B(4) and A(4);
sig_137 <= B(5) and A(4);
sig_138 <= B(6) and A(4);
sig_139 <= B(7) and A(4);
sig_160 <= sig_125 xor sig_136;
sig_161 <= sig_125 and sig_136;
sig_162 <= sig_160 and sig_118;
sig_163 <= sig_160 or sig_118;
sig_164 <= sig_161 or sig_162;
sig_165 <= sig_130 xor sig_137;
sig_166 <= sig_130 and sig_137;
sig_167 <= sig_165 and sig_126;
sig_168 <= sig_165 xor sig_126;
sig_169 <= sig_166 or sig_167;
sig_170 <= sig_96 xor sig_138;
sig_171 <= sig_96 and sig_138;
sig_172 <= sig_170 and sig_131;
sig_173 <= sig_170 xor sig_131;
sig_174 <= sig_171 or sig_172;
sig_177 <= B(2) and A(5);
sig_178 <= B(3) and A(5);
sig_179 <= B(4) and A(5);
sig_180 <= B(5) and A(5);
sig_181 <= B(6) and A(5);
sig_182 <= B(7) and A(5);
sig_196 <= sig_162 xor sig_117;
sig_198 <= sig_163 xor sig_178;
sig_199 <= sig_163 and sig_178;
sig_200 <= sig_198 and sig_113;
sig_201 <= sig_198 xor sig_113;
sig_202 <= sig_199 or sig_200;
sig_203 <= sig_168 xor sig_179;
sig_204 <= sig_168 and sig_179;
sig_205 <= sig_203 and sig_164;
sig_206 <= sig_203 xor sig_164;
sig_207 <= sig_204 or sig_205;
sig_208 <= sig_173 xor sig_180;
sig_209 <= sig_173 and sig_180;
sig_210 <= sig_208 and sig_169;
sig_211 <= sig_208 xor sig_169;
sig_212 <= sig_209 or sig_210;
sig_213 <= sig_139 xor sig_181;
sig_214 <= sig_139 and sig_181;
sig_215 <= sig_213 and sig_174;
sig_216 <= sig_213 xor sig_174;
sig_217 <= sig_214 or sig_215;
sig_219 <= B(1) and A(6);
sig_220 <= B(2) and A(6);
sig_221 <= B(3) and A(6);
sig_222 <= B(4) and A(6);
sig_223 <= B(5) and A(6);
sig_224 <= B(6) and A(6);
sig_225 <= B(7) and A(6);
sig_231 <= sig_196 xor sig_219;
sig_232 <= sig_196 and sig_219;
sig_236 <= sig_201 xor sig_220;
sig_237 <= sig_201 and sig_220;
sig_238 <= sig_236 and sig_177;
sig_239 <= sig_236 xor sig_177;
sig_240 <= sig_237 or sig_238;
sig_241 <= sig_206 xor sig_221;
sig_242 <= sig_206 and sig_221;
sig_243 <= sig_241 and sig_202;
sig_244 <= sig_241 xor sig_202;
sig_245 <= sig_242 or sig_243;
sig_246 <= sig_211 xor sig_222;
sig_247 <= sig_211 and sig_222;
sig_248 <= sig_246 and sig_207;
sig_249 <= sig_246 xor sig_207;
sig_250 <= sig_247 or sig_248;
sig_251 <= sig_216 xor sig_223;
sig_252 <= sig_216 and sig_223;
sig_253 <= sig_251 and sig_212;
sig_254 <= sig_251 xor sig_212;
sig_255 <= sig_252 or sig_253;
sig_256 <= sig_182 xor sig_224;
sig_257 <= sig_182 and sig_224;
sig_258 <= sig_256 and sig_217;
sig_259 <= sig_256 xor sig_217;
sig_260 <= sig_257 or sig_258;
sig_261 <= B(0) and A(7);
sig_262 <= B(1) and A(7);
sig_263 <= B(2) and A(7);
sig_264 <= B(3) and A(7);
sig_265 <= B(4) and A(7);
sig_266 <= B(5) and A(7);
sig_267 <= B(6) and A(7);
sig_268 <= B(7) and A(7);
sig_273 <= sig_225 and sig_267;
sig_274 <= sig_239 xor sig_262;
sig_275 <= sig_239 and sig_262;
sig_276 <= sig_274 and sig_232;
sig_277 <= sig_274 or sig_232;
sig_278 <= sig_275 or sig_276;
sig_279 <= sig_244 xor sig_263;
sig_280 <= sig_244 and sig_263;
sig_281 <= sig_279 and sig_240;
sig_282 <= sig_279 xor sig_240;
sig_283 <= sig_280 or sig_281;
sig_284 <= sig_249 xor sig_264;
sig_285 <= sig_249 and sig_264;
sig_286 <= sig_284 and sig_245;
sig_287 <= sig_284 xor sig_245;
sig_288 <= sig_285 or sig_286;
sig_289 <= sig_254 xor sig_265;
sig_290 <= sig_254 and sig_265;
sig_291 <= sig_289 and sig_250;
sig_292 <= sig_289 xor sig_250;
sig_293 <= sig_290 or sig_291;
sig_294 <= sig_259 xor sig_266;
sig_295 <= sig_259 and sig_266;
sig_296 <= sig_294 and sig_255;
sig_297 <= sig_294 xor sig_255;
sig_298 <= sig_295 or sig_296;
sig_299 <= sig_225 xor sig_267;
sig_301 <= sig_299 and sig_260;
sig_302 <= sig_299 xor sig_260;
sig_303 <= sig_273 or sig_301;
sig_306 <= sig_282 xor sig_278;
sig_307 <= sig_282 and sig_278;
sig_311 <= sig_287 xor sig_283;
sig_312 <= sig_287 and sig_283;
sig_313 <= sig_311 and sig_307;
sig_314 <= sig_311 xor sig_307;
sig_315 <= sig_312 or sig_313;
sig_316 <= sig_292 xor sig_288;
sig_317 <= sig_292 and sig_288;
sig_318 <= sig_316 and sig_315;
sig_319 <= sig_316 xor sig_315;
sig_320 <= sig_317 or sig_318;
sig_321 <= sig_297 xor sig_293;
sig_322 <= sig_297 and sig_293;
sig_323 <= sig_321 and sig_320;
sig_324 <= sig_321 xor sig_320;
sig_325 <= sig_322 or sig_323;
sig_326 <= sig_302 xor sig_298;
sig_327 <= sig_302 and sig_298;
sig_328 <= sig_326 and sig_325;
sig_329 <= sig_326 xor sig_325;
sig_330 <= sig_327 or sig_328;
sig_331 <= sig_268 xor sig_303;
sig_332 <= A(7) and sig_303;
sig_333 <= sig_268 and sig_330;
sig_334 <= sig_331 xor sig_330;
sig_335 <= sig_332 or sig_333;
O(15) <= sig_335;
O(14) <= sig_334;
O(13) <= sig_329;
O(12) <= sig_324;
O(11) <= sig_319;
O(10) <= sig_314;
O(9) <= sig_306;
O(8) <= sig_277;
O(7) <= sig_261;
O(6) <= sig_231;
O(5) <= sig_199;
O(4) <= sig_264;
O(3) <= sig_117;
O(2) <= sig_260;
O(1) <= sig_163;
O(0) <= sig_177;
end mul8u_197B_struct;
