entity mul8u_LK8 is
port (A : in std_logic_vector (7 downto 0);
B : in std_logic_vector (7 downto 0);
O : out std_logic_vector (15 downto 0)
);
end mul8u_LK8;
architecture mul8u_LK8_struct of mul8u_LK8 is
signal sig_19,sig_20,sig_21,sig_22,sig_23,sig_26,sig_27,sig_28,sig_29,sig_30,sig_31,sig_35,sig_36,sig_37,sig_38,sig_39,sig_40,sig_41,sig_42,sig_43: std_logic;
signal sig_44,sig_45,sig_47,sig_48,sig_49,sig_50,sig_51,sig_52,sig_53,sig_59,sig_60,sig_64,sig_65,sig_66,sig_67,sig_68,sig_69,sig_70,sig_71,sig_72: std_logic;
signal sig_73,sig_74,sig_75,sig_76,sig_77,sig_78,sig_79,sig_80,sig_81,sig_82,sig_83,sig_84,sig_85,sig_87,sig_88,sig_89,sig_90,sig_91,sig_92,sig_93: std_logic;
signal sig_94,sig_95,sig_96,sig_97,sig_98,sig_102,sig_103,sig_104,sig_105,sig_106,sig_107,sig_108,sig_109,sig_110,sig_111,sig_112,sig_113,sig_114,sig_115,sig_116: std_logic;
signal sig_117,sig_118,sig_119,sig_120,sig_121,sig_122,sig_123,sig_124,sig_125,sig_126,sig_127,sig_128,sig_129,sig_130,sig_131,sig_132,sig_133,sig_134,sig_135,sig_136: std_logic;
signal sig_137,sig_138,sig_139,sig_140,sig_141,sig_142,sig_143,sig_144,sig_145,sig_146,sig_147,sig_148,sig_149,sig_150,sig_151,sig_152,sig_153,sig_154,sig_155,sig_156: std_logic;
signal sig_157,sig_158,sig_159,sig_160,sig_161,sig_162,sig_163,sig_164,sig_165,sig_166,sig_167,sig_168,sig_169,sig_170,sig_171,sig_172,sig_173,sig_174,sig_175,sig_176: std_logic;
signal sig_177,sig_178,sig_179,sig_180,sig_181,sig_182,sig_183,sig_184,sig_185,sig_186,sig_187,sig_188,sig_189,sig_190,sig_191,sig_192,sig_193,sig_194,sig_195,sig_196: std_logic;
signal sig_197,sig_198,sig_199,sig_200,sig_201,sig_202,sig_203,sig_204,sig_205,sig_206,sig_207,sig_208,sig_209,sig_210,sig_211,sig_212,sig_213,sig_214,sig_215,sig_216: std_logic;
signal sig_217,sig_218,sig_219,sig_220,sig_221,sig_222,sig_223,sig_224,sig_225,sig_226,sig_227,sig_228,sig_229,sig_230,sig_231,sig_232,sig_233,sig_234,sig_235,sig_236: std_logic;
signal sig_237,sig_238,sig_239,sig_240,sig_241,sig_242,sig_243,sig_244,sig_245,sig_246,sig_247,sig_248,sig_249,sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256: std_logic;
signal sig_257,sig_258,sig_259,sig_260,sig_261,sig_262,sig_263,sig_264,sig_265,sig_266,sig_267,sig_268,sig_269,sig_270,sig_271,sig_272,sig_273,sig_274,sig_275,sig_276: std_logic;
signal sig_277,sig_278,sig_279,sig_280,sig_281,sig_282,sig_283,sig_284,sig_285,sig_286,sig_287,sig_288,sig_289,sig_290,sig_291,sig_292,sig_293,sig_294,sig_295,sig_296: std_logic;
signal sig_297,sig_298,sig_299,sig_300,sig_301,sig_302,sig_303,sig_304,sig_305,sig_306,sig_307,sig_308,sig_309,sig_310,sig_311,sig_312,sig_313,sig_314,sig_315,sig_316: std_logic;
signal sig_317,sig_318,sig_319,sig_320,sig_321,sig_322,sig_323,sig_324,sig_325,sig_326,sig_327,sig_328,sig_329,sig_330,sig_331,sig_332,sig_333,sig_334,sig_335: std_logic;
begin
sig_19 <= B(3) and A(0);
sig_20 <= B(4) and A(0);
sig_21 <= B(5) and A(0);
sig_22 <= B(6) and A(0);
sig_23 <= B(7) and A(0);
sig_26 <= B(2) and A(1);
sig_27 <= B(3) and A(1);
sig_28 <= B(4) and A(1);
sig_29 <= B(5) and A(1);
sig_30 <= B(6) and A(1);
sig_31 <= B(7) and A(1);
sig_35 <= B(6) and sig_31;
sig_36 <= sig_19 or sig_26;
sig_37 <= sig_19 and sig_26;
sig_38 <= sig_20 xor sig_27;
sig_39 <= sig_20 and sig_27;
sig_40 <= sig_21 xor sig_28;
sig_41 <= sig_21 and sig_28;
sig_42 <= sig_22 xor sig_29;
sig_43 <= sig_22 and sig_29;
sig_44 <= sig_23 xor sig_30;
sig_45 <= A(0) and sig_35;
sig_47 <= B(1) and A(2);
sig_48 <= B(2) and A(2);
sig_49 <= B(3) and A(2);
sig_50 <= B(4) and A(2);
sig_51 <= B(5) and A(2);
sig_52 <= B(6) and A(2);
sig_53 <= B(7) and A(2);
sig_59 <= sig_36 or sig_47;
sig_60 <= sig_36 and sig_47;
sig_64 <= sig_38 xor sig_48;
sig_65 <= sig_38 and sig_48;
sig_66 <= sig_64 and sig_37;
sig_67 <= sig_64 xor sig_37;
sig_68 <= sig_65 or sig_66;
sig_69 <= sig_40 xor sig_49;
sig_70 <= sig_40 and sig_49;
sig_71 <= sig_69 and sig_39;
sig_72 <= sig_69 xor sig_39;
sig_73 <= sig_70 or sig_71;
sig_74 <= sig_42 xor sig_50;
sig_75 <= sig_42 and sig_50;
sig_76 <= sig_74 and sig_41;
sig_77 <= sig_74 xor sig_41;
sig_78 <= sig_75 or sig_76;
sig_79 <= sig_44 xor sig_51;
sig_80 <= sig_44 and sig_51;
sig_81 <= sig_79 and sig_43;
sig_82 <= sig_79 xor sig_43;
sig_83 <= sig_80 or sig_81;
sig_84 <= sig_31 xor sig_52;
sig_85 <= sig_35 and sig_52;
sig_87 <= sig_84 xor sig_45;
sig_88 <= sig_85 or sig_45;
sig_89 <= B(0) and A(3);
sig_90 <= B(1) and A(3);
sig_91 <= B(2) and A(3);
sig_92 <= B(3) and A(3);
sig_93 <= B(4) and A(3);
sig_94 <= B(5) and A(3);
sig_95 <= B(6) and A(3);
sig_96 <= B(7) and A(3);
sig_97 <= sig_59 or sig_89;
sig_98 <= sig_59 and sig_89;
sig_102 <= sig_67 xor sig_90;
sig_103 <= sig_67 and sig_90;
sig_104 <= sig_102 and sig_60;
sig_105 <= sig_102 xor sig_60;
sig_106 <= sig_103 or sig_104;
sig_107 <= sig_72 xor sig_91;
sig_108 <= sig_72 and sig_91;
sig_109 <= sig_107 and sig_68;
sig_110 <= sig_107 xor sig_68;
sig_111 <= sig_108 or sig_109;
sig_112 <= sig_77 xor sig_92;
sig_113 <= sig_77 and sig_92;
sig_114 <= sig_112 and sig_73;
sig_115 <= sig_112 xor sig_73;
sig_116 <= sig_113 or sig_114;
sig_117 <= sig_82 xor sig_93;
sig_118 <= sig_82 and sig_93;
sig_119 <= sig_117 and sig_78;
sig_120 <= sig_117 xor sig_78;
sig_121 <= sig_118 or sig_119;
sig_122 <= sig_87 xor sig_94;
sig_123 <= sig_87 and sig_94;
sig_124 <= sig_122 and sig_83;
sig_125 <= sig_122 xor sig_83;
sig_126 <= sig_123 or sig_124;
sig_127 <= sig_53 xor sig_95;
sig_128 <= sig_53 and sig_95;
sig_129 <= sig_127 and sig_88;
sig_130 <= sig_127 xor sig_88;
sig_131 <= sig_128 or sig_129;
sig_132 <= B(0) and A(4);
sig_133 <= B(1) and A(4);
sig_134 <= B(2) and A(4);
sig_135 <= B(3) and A(4);
sig_136 <= B(4) and A(4);
sig_137 <= B(5) and A(4);
sig_138 <= B(6) and A(4);
sig_139 <= B(7) and A(4);
sig_140 <= sig_105 xor sig_132;
sig_141 <= sig_105 and sig_132;
sig_142 <= sig_140 and sig_98;
sig_143 <= sig_140 xor sig_98;
sig_144 <= sig_141 or sig_142;
sig_145 <= sig_110 xor sig_133;
sig_146 <= sig_110 and sig_133;
sig_147 <= sig_145 and sig_106;
sig_148 <= sig_145 xor sig_106;
sig_149 <= sig_146 or sig_147;
sig_150 <= sig_115 xor sig_134;
sig_151 <= sig_115 and sig_134;
sig_152 <= sig_150 and sig_111;
sig_153 <= sig_150 xor sig_111;
sig_154 <= sig_151 or sig_152;
sig_155 <= sig_120 xor sig_135;
sig_156 <= sig_120 and sig_135;
sig_157 <= sig_155 and sig_116;
sig_158 <= sig_155 xor sig_116;
sig_159 <= sig_156 or sig_157;
sig_160 <= sig_125 xor sig_136;
sig_161 <= sig_125 and sig_136;
sig_162 <= sig_160 and sig_121;
sig_163 <= sig_160 xor sig_121;
sig_164 <= sig_161 or sig_162;
sig_165 <= sig_130 xor sig_137;
sig_166 <= sig_130 and sig_137;
sig_167 <= sig_165 and sig_126;
sig_168 <= sig_165 xor sig_126;
sig_169 <= sig_166 or sig_167;
sig_170 <= sig_96 xor sig_138;
sig_171 <= sig_96 and sig_138;
sig_172 <= sig_170 and sig_131;
sig_173 <= sig_170 xor sig_131;
sig_174 <= sig_171 or sig_172;
sig_175 <= B(0) and A(5);
sig_176 <= B(1) and A(5);
sig_177 <= B(2) and A(5);
sig_178 <= B(3) and A(5);
sig_179 <= B(4) and A(5);
sig_180 <= B(5) and A(5);
sig_181 <= B(6) and A(5);
sig_182 <= B(7) and A(5);
sig_183 <= sig_148 xor sig_175;
sig_184 <= sig_148 and sig_175;
sig_185 <= sig_183 and sig_144;
sig_186 <= sig_183 xor sig_144;
sig_187 <= sig_184 or sig_185;
sig_188 <= sig_153 xor sig_176;
sig_189 <= sig_153 and sig_176;
sig_190 <= sig_188 and sig_149;
sig_191 <= sig_188 xor sig_149;
sig_192 <= sig_189 or sig_190;
sig_193 <= sig_158 xor sig_177;
sig_194 <= sig_158 and sig_177;
sig_195 <= sig_193 and sig_154;
sig_196 <= sig_193 xor sig_154;
sig_197 <= sig_194 or sig_195;
sig_198 <= sig_163 xor sig_178;
sig_199 <= sig_163 and sig_178;
sig_200 <= sig_198 and sig_159;
sig_201 <= sig_198 xor sig_159;
sig_202 <= sig_199 or sig_200;
sig_203 <= sig_168 xor sig_179;
sig_204 <= sig_168 and sig_179;
sig_205 <= sig_203 and sig_164;
sig_206 <= sig_203 xor sig_164;
sig_207 <= sig_204 or sig_205;
sig_208 <= sig_173 xor sig_180;
sig_209 <= sig_173 and sig_180;
sig_210 <= sig_208 and sig_169;
sig_211 <= sig_208 xor sig_169;
sig_212 <= sig_209 or sig_210;
sig_213 <= sig_139 xor sig_181;
sig_214 <= sig_139 and sig_181;
sig_215 <= sig_213 and sig_174;
sig_216 <= sig_213 xor sig_174;
sig_217 <= sig_214 or sig_215;
sig_218 <= B(0) and A(6);
sig_219 <= B(1) and A(6);
sig_220 <= B(2) and A(6);
sig_221 <= B(3) and A(6);
sig_222 <= B(4) and A(6);
sig_223 <= B(5) and A(6);
sig_224 <= B(6) and A(6);
sig_225 <= B(7) and A(6);
sig_226 <= sig_191 xor sig_218;
sig_227 <= sig_191 and sig_218;
sig_228 <= sig_226 and sig_187;
sig_229 <= sig_226 xor sig_187;
sig_230 <= sig_227 or sig_228;
sig_231 <= sig_196 xor sig_219;
sig_232 <= sig_196 and sig_219;
sig_233 <= sig_231 and sig_192;
sig_234 <= sig_231 xor sig_192;
sig_235 <= sig_232 or sig_233;
sig_236 <= sig_201 xor sig_220;
sig_237 <= sig_201 and sig_220;
sig_238 <= sig_236 and sig_197;
sig_239 <= sig_236 xor sig_197;
sig_240 <= sig_237 or sig_238;
sig_241 <= sig_206 xor sig_221;
sig_242 <= sig_206 and sig_221;
sig_243 <= sig_241 and sig_202;
sig_244 <= sig_241 xor sig_202;
sig_245 <= sig_242 or sig_243;
sig_246 <= sig_211 xor sig_222;
sig_247 <= sig_211 and sig_222;
sig_248 <= sig_246 and sig_207;
sig_249 <= sig_246 xor sig_207;
sig_250 <= sig_247 or sig_248;
sig_251 <= sig_216 xor sig_223;
sig_252 <= sig_216 and sig_223;
sig_253 <= sig_251 and sig_212;
sig_254 <= sig_251 xor sig_212;
sig_255 <= sig_252 or sig_253;
sig_256 <= sig_182 xor sig_224;
sig_257 <= sig_182 and sig_224;
sig_258 <= sig_256 and sig_217;
sig_259 <= sig_256 xor sig_217;
sig_260 <= sig_257 or sig_258;
sig_261 <= B(0) and A(7);
sig_262 <= B(1) and A(7);
sig_263 <= B(2) and A(7);
sig_264 <= B(3) and A(7);
sig_265 <= B(4) and A(7);
sig_266 <= B(5) and A(7);
sig_267 <= B(6) and A(7);
sig_268 <= B(7) and A(7);
sig_269 <= sig_234 xor sig_261;
sig_270 <= sig_234 and sig_261;
sig_271 <= sig_269 and sig_230;
sig_272 <= sig_269 xor sig_230;
sig_273 <= sig_270 or sig_271;
sig_274 <= sig_239 xor sig_262;
sig_275 <= sig_239 and sig_262;
sig_276 <= sig_274 and sig_235;
sig_277 <= sig_274 xor sig_235;
sig_278 <= sig_275 or sig_276;
sig_279 <= sig_244 xor sig_263;
sig_280 <= sig_244 and sig_263;
sig_281 <= sig_279 and sig_240;
sig_282 <= sig_279 xor sig_240;
sig_283 <= sig_280 or sig_281;
sig_284 <= sig_249 xor sig_264;
sig_285 <= sig_249 and sig_264;
sig_286 <= sig_284 and sig_245;
sig_287 <= sig_284 xor sig_245;
sig_288 <= sig_285 or sig_286;
sig_289 <= sig_254 xor sig_265;
sig_290 <= sig_254 and sig_265;
sig_291 <= sig_289 and sig_250;
sig_292 <= sig_289 xor sig_250;
sig_293 <= sig_290 or sig_291;
sig_294 <= sig_259 xor sig_266;
sig_295 <= sig_259 and sig_266;
sig_296 <= sig_294 and sig_255;
sig_297 <= sig_294 xor sig_255;
sig_298 <= sig_295 or sig_296;
sig_299 <= sig_225 xor sig_267;
sig_300 <= sig_225 and sig_267;
sig_301 <= sig_299 and sig_260;
sig_302 <= sig_299 xor sig_260;
sig_303 <= sig_300 or sig_301;
sig_304 <= sig_277 xor sig_273;
sig_305 <= sig_277 and sig_273;
sig_306 <= sig_282 xor sig_278;
sig_307 <= sig_282 and sig_278;
sig_308 <= sig_306 and sig_305;
sig_309 <= sig_306 xor sig_305;
sig_310 <= sig_307 or sig_308;
sig_311 <= sig_287 xor sig_283;
sig_312 <= sig_287 and sig_283;
sig_313 <= sig_311 and sig_310;
sig_314 <= sig_311 xor sig_310;
sig_315 <= sig_312 or sig_313;
sig_316 <= sig_292 xor sig_288;
sig_317 <= sig_292 and sig_288;
sig_318 <= sig_316 and sig_315;
sig_319 <= sig_316 xor sig_315;
sig_320 <= sig_317 or sig_318;
sig_321 <= sig_297 xor sig_293;
sig_322 <= sig_297 and sig_293;
sig_323 <= sig_321 and sig_320;
sig_324 <= sig_321 xor sig_320;
sig_325 <= sig_322 or sig_323;
sig_326 <= sig_302 xor sig_298;
sig_327 <= sig_302 and sig_298;
sig_328 <= sig_326 and sig_325;
sig_329 <= sig_326 xor sig_325;
sig_330 <= sig_327 or sig_328;
sig_331 <= sig_268 xor sig_303;
sig_332 <= A(7) and sig_303;
sig_333 <= sig_331 and sig_330;
sig_334 <= sig_331 xor sig_330;
sig_335 <= sig_332 or sig_333;
O(15) <= sig_335;
O(14) <= sig_334;
O(13) <= sig_329;
O(12) <= sig_324;
O(11) <= sig_319;
O(10) <= sig_314;
O(9) <= sig_309;
O(8) <= sig_304;
O(7) <= sig_272;
O(6) <= sig_229;
O(5) <= sig_186;
O(4) <= sig_143;
O(3) <= sig_97;
O(2) <= 1'b0;
O(1) <= sig_97;
O(0) <= 1'b0;
end mul8u_LK8_struct;
